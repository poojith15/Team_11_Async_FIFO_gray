khvouvoyy
